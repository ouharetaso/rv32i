

module cpu (
    inout  b_membus[31:0],
    output o_memaddr[31:0]
);
    


endmodule